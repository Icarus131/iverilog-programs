module and1(input wire a,b,output wire x);
assign y = a&b;

endmodule
