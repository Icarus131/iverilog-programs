module and1(input wire c,b,output wire x);
assign x = c&b;

endmodule
