module not1(input wire a,output wire x);
assign x = ~a;

endmodule
