module xor1(input wire a,b,output wire x,y);
assign y = a^b;

endmodule
